`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 09.09.2023 15:53:24
// Design Name: 
// Module Name: lab2_assignment_multiplexer
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module lab2_assignment_multiplexer(
    input [5:0] DR,
    input [5:0] NR,
    input Button,
    output [5:0] Z
    );
endmodule
